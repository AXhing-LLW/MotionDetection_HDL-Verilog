// megafunction wizard: %Shift register (RAM-based)%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altshift_taps 

// ============================================================
// File Name: Tap_1.v
// Megafunction Name(s):
// 			altshift_taps
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 5.1 Build 213 01/19/2006 SP 1 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2006 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module Tap_1 (
	clken,
	clock,
	shiftin,
	shiftout,
	taps);

	input	  clken;
	input	  clock;
	input	  shiftin;
	output	  shiftout;
	output	[10:0]  taps;

	wire [10:0] sub_wire0;
	wire [0:0] sub_wire1;
	wire [10:0] taps = sub_wire0[10:0];
	wire [0:0] sub_wire2 = sub_wire1[0:0];
	wire  shiftout = sub_wire2;
	wire  sub_wire3 = shiftin;
	wire  sub_wire4 = sub_wire3;

	altshift_taps	altshift_taps_component (
				.clken (clken),
				.clock (clock),
				.shiftin (sub_wire4),
				.taps (sub_wire0),
				.shiftout (sub_wire1));
	defparam
		altshift_taps_component.lpm_type = "altshift_taps",
		altshift_taps_component.number_of_taps = 11,
		altshift_taps_component.tap_distance = 640,
		altshift_taps_component.width = 1;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: CLKEN NUMERIC "1"
// Retrieval info: PRIVATE: GROUP_TAPS NUMERIC "0"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
// Retrieval info: PRIVATE: NUMBER_OF_TAPS NUMERIC "11"
// Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "0"
// Retrieval info: PRIVATE: TAP_DISTANCE NUMERIC "640"
// Retrieval info: PRIVATE: WIDTH NUMERIC "1"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altshift_taps"
// Retrieval info: CONSTANT: NUMBER_OF_TAPS NUMERIC "11"
// Retrieval info: CONSTANT: TAP_DISTANCE NUMERIC "640"
// Retrieval info: CONSTANT: WIDTH NUMERIC "1"
// Retrieval info: USED_PORT: clken 0 0 0 0 INPUT VCC clken
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL clock
// Retrieval info: USED_PORT: shiftin 0 0 0 0 INPUT NODEFVAL shiftin
// Retrieval info: USED_PORT: shiftout 0 0 0 0 OUTPUT NODEFVAL shiftout
// Retrieval info: USED_PORT: taps 0 0 11 0 OUTPUT NODEFVAL taps[10..0]
// Retrieval info: CONNECT: @shiftin 0 0 1 0 shiftin 0 0 0 0
// Retrieval info: CONNECT: shiftout 0 0 0 0 @shiftout 0 0 1 0
// Retrieval info: CONNECT: taps 0 0 11 0 @taps 0 0 11 0
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: CONNECT: @clken 0 0 0 0 clken 0 0 0 0
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: GEN_FILE: TYPE_NORMAL Tap_1.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL Tap_1.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL Tap_1.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL Tap_1.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL Tap_1_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL Tap_1_bb.v FALSE
